LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;

ENTITY TEST_TB IS
END TEST_TB;

ARCHITECTURE TRY OF TEST_TB IS
	COMPONENT TEST
		PORT( 
			CLK, CLR, ES: IN STD_LOGIC;
			D: IN STD_LOGIC_VECTOR(6 DOWNTO 0);
			OP: IN STD_LOGIC_VECTOR(1 DOWNTO 0);
			Q: INOUT STD_LOGIC_VECTOR(6 DOWNTO 0)
		);
	END COMPONENT;

	SIGNAL CLK, CLR, ES : STD_LOGIC;
	SIGNAL D : STD_LOGIC_VECTOR(6 DOWNTO 0);
	SIGNAL OP : STD_LOGIC_VECTOR(1 DOWNTO 0);
	SIGNAL Q : STD_LOGIC_VECTOR(6 DOWNTO 0);

	SIGNAL CLK_PERIOD : time := 10ns; -- Reloj de 100MHz

	BEGIN
		REGISTRO : TEST PORT MAP (CLK => CLK, CLR => CLR, ES => ES, D => D, OP => OP, Q => Q);

		PROCESS
			BEGIN
				CLK <= '0';
				WAIT FOR 5 NS;
				CLK <= '1';
				WAIT FOR 5 NS;
		END PROCESS;

		PROCESS
			BEGIN
				ES <= '1';
				WAIT FOR 3 NS;
				ES <= '0';
				WAIT FOR 3 NS;
		END PROCESS;

		PROCESS
			BEGIN
				OP <= "00";
				WAIT FOR 4 NS;
				OP <= "01";
				WAIT FOR 4 NS;
				OP <= "10";
				WAIT FOR 4 NS;
				OP <= "11";
				WAIT FOR 4 NS;
		END PROCESS;

		PROCESS
			BEGIN
				D <= "1011001";
				WAIT FOR 7 NS;
				D <= "0010110";
				WAIT FOR 7 NS;
		END PROCESS;

		-- ASSERT FALSE REPORT "REACHED END OF TEST";
END TRY;