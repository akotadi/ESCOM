LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.ALL;

-- INCLUIR PAQUETE CON CONSTANTES DE OPCODE, FUNCODE Y REGISTROS
LIBRARY WORK;
USE WORK.PKG_ESCOMIPS.ALL;

ENTITY CONTROL IS
	GENERIC( 
		BC : INTEGER := 20;
		ADR_F : INTEGER := 4;
		ADR_OP : INTEGER := 5
	);

	Port ( 
		FUNCODE : IN STD_LOGIC_VECTOR (ADR_F-1 DOWNTO 0);
		OPCODE : IN STD_LOGIC_VECTOR (ADR_OP-1 DOWNTO 0);
		Z, C, N, OV : IN STD_LOGIC;
		LF, CLK, CLR : IN STD_LOGIC;
		BCTRL : OUT STD_LOGIC_VECTOR (BC-1 DOWNTO 0)
	);
END CONTROL;

ARCHITECTURE UNIDAD OF CONTROL IS

-- UNIDAD DE CONTROL
TYPE ESTADOS IS ( A );
SIGNAL EDO_ACT, EDO_SGTE : ESTADOS;
-- MEMORIA DE MICROCÓDIGO DE FUNCIÓN
TYPE MEM_FUNCT IS ARRAY( 0 TO (2**ARD_F)-1 ) OF STD_LOGIC_VECTOR( BCTRL'RANGE );
CONSTANT MICRO_COD_FU : MEM_FUNCT := (
	-- COPIAR DEL DOCUMENTO
	"00000100110000011001"; -- ADD
	"00000100110000111001"; -- SUB
	"00000100110000000001"; -- AND
	"00000100110000001001"; -- OR
	"00000100110000010001"; -- XOR
	"00000100110001101001"; -- NAND
	"00000100110001100001"; -- NOR
	"00000100110001010001"; -- XNOR
	"00000100110001101001"; -- NOT
	"00000011000000000000"; -- SLL
	"00000010000000000000"; -- SRL
	OTHERS => ( OTHERS => '0' )
);
-- MEMORIA DE MICROCÓDIGO DE OPERACIÓN
TYPE MEM_OPT IS ARRAY( 0 TO (2**ARD_OP)-1 ) OF STD_LOGIC_VECTOR( BCTRL'RANGE );
CONSTANT MICRO_COD_OPT : MEM_OPT := (
	"00001000010000111000"; -- Bcond
	"00000000100000000000"; -- LI
	"00000100100000000100"; -- LWI
	"00001000000000000110"; -- SWI
	"00001000001010011010"; -- SW
	"00000100110010011001"; -- ADDI
	"00000100110010111001"; -- SUBI
	"00000100111010000001"; -- ANDI
	"00000100111010001001"; -- ORI
	"00000100111010010001"; -- XORI
	"00000100111011101001"; -- NANDI
	"00000100111011100001"; -- NORI
	"00000100111011010001"; -- XNORI
	"00110000000110011001"; -- BEQI
	"00110000000110011001"; -- BNEI
	"00110000000110011001"; -- BLTI
	"00110000000110011001"; -- BLETI
	"00110000000110011001"; -- BGTI
	"00110000000110011001"; -- BGETI
	"00100000000000000000"; -- B
	"10100000000000000000"; -- CALL
	"01000000000000000000"; -- RET
	"00000000000000000000"; -- NOP 
	"00000100011010011000"; -- LW
	OTHERS => ( OTHERS => '0' )
);
-- SEÑALES DEL DECODIFICADOR DE INSTRUCCIÓN
SIGNAL TIPOR, BEQI, BNEQI, BLTI, BLETI, BGTI, BGETI : STD_LOGIC;
-- SEÑALES DEL REGISTRO DE ESTADO
SIGNAL RZ, RC, RN, ROV : STD_LOGIC;
-- SEÑALES DE CONDICIÓN
SIGNAL EQ, NEQ, LTI, LETI, GTI, GETI : STD_LOGIC;
-- SEÑALES DE UNIDAD DE CONTROL
SIGNAL SDOPC, SM : STD_LOGIC;
-- SEÑAL DE MICROCÓDIGO DE FUNCIÓN
SIGNAL DF : STD_LOGIC_VECTOR( BCTRL'RANGE );
-- SEÑAL DE MICROCÓDIGO DE OPERACIÓN
SIGNAL S_OPCODE : STD_LOGIC_VECTOR( OPCODE'RANGE );
SIGNAL D : STD_LOGIC_VECTOR( BCTRL'RANGE );


-- MOVER A PAQUETE JUNTO CON LOS DEMÁS CÓDIGOS 
CONSTANT OPCODE_BEQI : STD_LOGIC_VECTOR( 4 DOWNTO 0 ) := "01101";
CONSTANT OPCODE_BNEQI : STD_LOGIC_VECTOR( 4 DOWNTO 0 ) := "01110";
CONSTANT OPCODE_BLTI : STD_LOGIC_VECTOR( 4 DOWNTO 0 ) := "01111";
CONSTANT OPCODE_BLETI : STD_LOGIC_VECTOR( 4 DOWNTO 0 ) := "10000";
CONSTANT OPCODE_BGTI : STD_LOGIC_VECTOR( 4 DOWNTO 0 ) := "10001";
CONSTANT OPCODE_BGETI : STD_LOGIC_VECTOR( 4 DOWNTO 0 ) := "10010";

	BEGIN

		DF <= MICRO_COD_FU( CONV_INTEGER(FUN_CODE) );

		S_OPCODE <= OPCODE WHEN ( SDOPC = '1' ) ELSE ( OTHERS => '0' ):
		D <= MICRO_COD_OPT( CONV_INTEGER(S_OPCODE) );

		BCTRL <= DF WHEN ( SM = '0' ) ELSE D;

		-- DECODIFICADOR DE INSTRUCCIÓN
		TIPOR <= '1' WHEN ( OPCODE = OPCODE_TIPOR ) ELSE '0';
		BEQI <= '1' WHEN ( OPCODE = OPCODE_BEQI ) ELSE '0';
		BNEQI <= '1' WHEN ( OPCODE = OPCODE_BNEQI ) ELSE '0';
		BLTI <= '1' WHEN ( OPCODE = OPCODE_BLTI ) ELSE '0';
		BLETI <= '1' WHEN ( OPCODE = OPCODE_BLETI ) ELSE '0';
		BGTI <= '1' WHEN ( OPCODE = OPCODE_BGTI ) ELSE '0';
		BGETI <= '1' WHEN ( OPCODE = OPCODE_BGETI ) ELSE '0';

		-- REGISTRO DE ESTADO
		PFLAGS : PROCESS ( CLK, CLR )
		BEGIN
			IF ( CLR = '1' ) THEN
				RZ <= '0';
				RC <= '0';
				RN <= '0';
				ROV <= '0';
			ELSIF ( FALLING_EDGE(CLK) ) THEN
				IF ( LF = '1' ) THEN
					RZ <= Z;
					RC <= C;
					RN <= N;
					ROV <= OV;
				END IF;
			END IF;
		END PROCESS PFLAGS;

		-- BLOQUE DE CONDICIÓN
		EQ <= RZ;
		NEQ <= NOT RZ;
		LTI <= ( NOT RZ ) AND ( RN XOR ROV );
		LETI <= RZ OR ( RN XOR ROV );
		GTI <= ( NOT RZ ) AND NOT ( RN XOR ROV);
		GETI <= RZ OR NOT ( RN XOR ROV);

		-- UNIDAD DE CONTROL

		TRANSICION : PROCESS ( CLK, CLR )
		BEGIN
			IF ( CLR = '1' ) THEN
				EDO_ACT <= A;
			ELSIF ( RISING_EDGE(CLK) ) THEN
				EDO_ACT <= EDO_SGTE;
			END IF;
		END PROCESS TRANSICION;

		AUTOMATA : PROCESS ( 
			TIPOR, BEQI, BNEQI, BLTI, BLETI, BGTI, BGETI, 
			EQ, NEQ, LTI, LETI, GTI, GETI 
		)
		BEGIN
			SM <= '0';
			SDOPC <= '0';
			CASE EDO_ACT IS
				WHEN A => 
					IF ( TIPOR = '1' ) THEN
						EDO_SGTE <= A;
					ELSE
						IF ( BEQI = '1' ) THEN
							IF ( CLK = '1' OR EQ = '0' ) THEN
								SM <= '1';
								EDO_SGTE <= A;
							ELSE 
								SM <= '1';
								SDOPC <= '1';
								EDO_SGTE <= A;
							END IF;
						ELSIF ( BNEQI = '1' ) THEN
							IF ( CLK = '1' OR NEQ = '0' ) THEN
								SM <= '1';
								EDO_SGTE <= A;
							ELSE 
								SM <= '1';
								SDOPC <= '1';
								EDO_SGTE <= A;
							END IF;
						ELSIF ( BLTI = '1' ) THEN
							IF ( CLK = '1' OR LTI = '0' ) THEN
								SM <= '1';
								EDO_SGTE <= A;
							ELSE 
								SM <= '1';
								SDOPC <= '1';
								EDO_SGTE <= A;
							END IF;
						ELSIF ( BLETI = '1' ) THEN
							IF ( CLK = '1' OR LETI = '0' ) THEN
								SM <= '1';
								EDO_SGTE <= A;
							ELSE 
								SM <= '1';
								SDOPC <= '1';
								EDO_SGTE <= A;
							END IF;
						ELSIF ( BGTI = '1' ) THEN
							IF ( CLK = '1' OR GTI = '0' ) THEN
								SM <= '1';
								EDO_SGTE <= A;
							ELSE 
								SM <= '1';
								SDOPC <= '1';
								EDO_SGTE <= A;
							END IF;
						ELSIF ( BGETI = '1' ) THEN
							IF ( CLK = '1' OR GETI = '0' ) THEN
								SM <= '1';
								EDO_SGTE <= A;
							ELSE 
								SM <= '1';
								SDOPC <= '1';
								EDO_SGTE <= A;
							END IF;
						ELSE
							SDOPC <= '1';
							SM <= '1';
							EDO_SGTE <= A;
						END IF;
					END IF;
			END CASE;
		END PROCESS AUTOMATA;

END UNIDAD;