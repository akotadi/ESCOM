LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.ALL;

ENTITY COMPUERTAS IS
	PORT(
			A:in STD_LOGIC;
			B:in STD_LOGIC;
			C:in STD_LOGIC;
			D:in STD_LOGIC;
			E:in STD_LOGIC;
			CAND: out STD_LOGIC;
			COR: out STD_LOGIC;
			CXOR: out STD_LOGIC;
			CNAND: out STD_LOGIC;
			CNOR: out STD_LOGIC;
			CXNOR: out STD_LOGIC
		);
END COMPUERTAS;

ARCHITECTURE BEHAVIORAL OF COMPUERTAS IS
	BEGIN
		CAND<= A AND B AND C AND D AND E;
		COR<= A OR B OR C OR D OR E;
		CXOR<= A XOR B XOR C XOR D XOR E;
		CNAND<= NOT CAND;
		CNOR<= NOT COR;
		CXNOR<= NOT CXOR;
	END BEHAVIORAL;