module compuertas ( 
	ams,
	bms,
	cinsc,
	cosc,
	cms,
	ssc,
	sms,
	amr,
	bmr,
	pirc,
	rmr,
	pmr,
	porc,
	rrc
	) ;

input  ams;
input  bms;
input  cinsc;
inout  cosc;
inout  cms;
inout  ssc;
inout  sms;
input  amr;
input  bmr;
input  pirc;
inout  rmr;
inout  pmr;
inout  porc;
inout  rrc;
