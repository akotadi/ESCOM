LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.ALL;

ENTITY COMPUERTAS IS
	PORT(
			A1: in STD_LOGIC;
			A2: in STD_LOGIC;
			A3: in STD_LOGIC;
			A4: in STD_LOGIC;
			B1: in STD_LOGIC;
			B2: in STD_LOGIC;
			B3: in STD_LOGIC;
			B4: in STD_LOGIC;
			Sel: in STD_LOGIC;
			Cout: out STD_LOGIC;
			S1: out STD_LOGIC;
			S2: out STD_LOGIC;
			S3: out STD_LOGIC;
			S4: out STD_LOGIC
			
		);

	ATTRIBUTE PIN_NUMBERS OF COMPUERTAS: ENTITY IS
	"A1:4 A2:3 A3:2 A4:1 B1:8 B2:7 B3:6 B4:5 Sel:9"
	& " S1:17 S2:16 S3:15 S4:14 Cout:18";
	


END COMPUERTAS;
ARCHITECTURE BEHAVIORAL OF COMPUERTAS IS
	BEGIN
		S1<= A1 XOR (B1 XOR Sel);
		S2<= (A2 XOR (B2 XOR Sel)) XOR Sel;
		S3<= (A3 XOR (B3 XOR Sel)) XOR Sel;
		S4<= (A4 XOR (B4 XOR Sel)) XOR Sel;
		Cout<= (((A4 XOR (B4 XOR Sel)) AND Sel) OR (A4 AND B4)) XOR Sel;
	END BEHAVIORAL;
