
LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;

ENTITY IMP_CRE IS
	PORT(
		CLK, CLR, EN : IN STD_LOGIC;
		Q : INOUT STD_LOGIC_VECTOR(9 DOWNTO 0)
	);

	ATTRIBUTE PIN_NUMBERS OF IMP_CRE : ENTITY IS 
		"CLK:1 "		&
		"EN:2 "			&
		"CLR:13 "		&
		"Q(0):15 "		&
		"Q(1):16 "		&
		"Q(2):17 "		&
		"Q(3):18 "		&
		"Q(4):19 "		&
		"Q(5):20 "		&
		"Q(6):21";
END IMP_CRE;

ARCHITECTURE PRACTICA OF IMP_CRE IS

	CONSTANT Symbol0 : STD_LOGIC_VECTOR(6 DOWNTO 0) := "0000001";
	CONSTANT Symbol1 : STD_LOGIC_VECTOR(6 DOWNTO 0) := "1001111";
	CONSTANT Symbol2 : STD_LOGIC_VECTOR(6 DOWNTO 0) := "0010010";
	CONSTANT Symbol3 : STD_LOGIC_VECTOR(6 DOWNTO 0) := "0000110";
	CONSTANT Symbol4 : STD_LOGIC_VECTOR(6 DOWNTO 0) := "1001100";
	CONSTANT Symbol5 : STD_LOGIC_VECTOR(6 DOWNTO 0) := "0100100";
	CONSTANT Symbol6 : STD_LOGIC_VECTOR(6 DOWNTO 0) := "0100000";
	CONSTANT Symbol7 : STD_LOGIC_VECTOR(6 DOWNTO 0) := "0001111";
	CONSTANT Symbol8 : STD_LOGIC_VECTOR(6 DOWNTO 0) := "0000000";
	CONSTANT Symbol9 : STD_LOGIC_VECTOR(6 DOWNTO 0) := "0000100";

	CONSTANT Label000 : STD_LOGIC_VECTOR(2 DOWNTO 0) := "000";
	CONSTANT Label001 : STD_LOGIC_VECTOR(2 DOWNTO 0) := "001";
	CONSTANT Label010 : STD_LOGIC_VECTOR(2 DOWNTO 0) := "010";
	CONSTANT Label011 : STD_LOGIC_VECTOR(2 DOWNTO 0) := "011";
	CONSTANT Label100 : STD_LOGIC_VECTOR(2 DOWNTO 0) := "100";
	CONSTANT Label101 : STD_LOGIC_VECTOR(2 DOWNTO 0) := "101";
	CONSTANT Label110 : STD_LOGIC_VECTOR(2 DOWNTO 0) := "110";
	CONSTANT Label111 : STD_LOGIC_VECTOR(2 DOWNTO 0) := "111";

	CONSTANT q0 : STD_LOGIC_VECTOR(9 DOWNTO 0) := Label000&Symbol2;
	CONSTANT q1 : STD_LOGIC_VECTOR(9 DOWNTO 0) := Label000&Symbol0;
	CONSTANT q2 : STD_LOGIC_VECTOR(9 DOWNTO 0) := Label000&Symbol1;
	CONSTANT q3 : STD_LOGIC_VECTOR(9 DOWNTO 0) := Label000&Symbol7;
	CONSTANT q4 : STD_LOGIC_VECTOR(9 DOWNTO 0) := Label000&Symbol6;
	CONSTANT q5 : STD_LOGIC_VECTOR(9 DOWNTO 0) := Label000&Symbol3;
	CONSTANT q6 : STD_LOGIC_VECTOR(9 DOWNTO 0) := Label001&Symbol0;
	CONSTANT q7 : STD_LOGIC_VECTOR(9 DOWNTO 0) := Label001&Symbol2;
	CONSTANT q8 : STD_LOGIC_VECTOR(9 DOWNTO 0) := Label010&Symbol0;
	CONSTANT q9 : STD_LOGIC_VECTOR(9 DOWNTO 0) := Label001&Symbol1;

	BEGIN

		PROCESS(CLK, CLR)
			BEGIN
				IF (CLR = '1') THEN
					Q <= q0;
				ELSIF RISING_EDGE(CLK) THEN
					IF ( EN = '1' ) THEN
						CASE Q IS
							WHEN q0 => Q <= q1;
							WHEN q1 => Q <= q2;
							WHEN q2 => Q <= q3;
							WHEN q3 => Q <= q4;
							WHEN q4 => Q <= q5;
							WHEN q5 => Q <= q6;
							WHEN q6 => Q <= q7;
							WHEN q7 => Q <= q8;
							WHEN q8 => Q <= q9;
							WHEN OTHERS => Q <= q0;
						END CASE;
					END IF;		
				END IF;
		END PROCESS;
END PRACTICA;