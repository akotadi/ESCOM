module compuertas ( 
	a,
	b,
	c,
	d,
	e,
	cand,
	cor,
	cxor,
	cnand,
	cnor,
	cxnor
	) ;

input  a;
input  b;
input  c;
input  d;
input  e;
inout  cand;
inout  cor;
inout  cxor;
inout  cnand;
inout  cnor;
inout  cxnor;
