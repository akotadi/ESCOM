LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.ALL;

ENTITY DETECTOR IS
	PORT(
		CLK, CLR, X: IN STD_LOGIC;
		AN: OUT STD_LOGIC;
		DISPLAY: OUT STD_LOGIC_VECTOR(6 DOWNTO 0)
	);

	ATTRIBUTE PIN_NUMBERS OF DETECTOR : ENTITY IS
		"CLK:1"			&
		"CLR:13"		&
		"X:11"			&
		"D(0):15"		&
		"D(1):16"		&
		"D(2):17"		&
		"D(3):18"		&
		"D(4):19"		&
		"D(5):20"		&
		"D(6):21"		&
		"AN:14";
END DETECTOR;

ARCHITECTURE PRACTICA OF DETECTOR IS

	SIGNAL Y, Qa, Qb : STD_LOGIC;

	CONSTANT SymbolA : STD_LOGIC_VECTOR(6 DOWNTO 0) := "0001000";
	CONSTANT SymbolE : STD_LOGIC_VECTOR(6 DOWNTO 0) := "0110000";

	BEGIN

		AN <= '0';

		PROCESS(CLK,CLR)
			BEGIN
				IF(CLR = '1') THEN
					Qa <= '0';
					Qb <= '0';
				ELSIF RISING_EDGE(CLK) THEN
					Qa <= ( NOT Qb AND X ) OR ( Qa AND X );
					Qb <= ( X AND Qa ) OR ( Qb AND Qa );
				END IF;
		END PROCESS;

		Y <= X AND ( NOT Qa ) AND Qb;

		DISPLAY <=
			SymbolA WHEN Y = '1' ELSE
			SymbolE;

END PRACTICA;