LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_UNSIGNED.ALL;

ENTITY ROM IS 

	GENERIC (
		BITS_BUS_DIR : INTEGER := 3;
		BITS_BUS_DATOS : INTEGER := 7
	);

	PORT(
		DIRECCION : IN STD_LOGIC_VECTOR( BITS_BUS_DIR-1 DOWNTO 0 );
		BUS_DATOS : OUT STD_LOGIC_VECTOR( BITS_BUS_DATOS-1 DOWNTO 0 );
		CS : IN STD_LOGIC
	);

END ROM;

ARCHITECTURE MEMORIA OF ROM IS 

	CONSTANT H : STD_LOGIC_VECTOR( 6 DOWNTO 0 ) := "1001000"; -- H
	CONSTANT O : STD_LOGIC_VECTOR( 6 DOWNTO 0 ) := "0000001"; -- O
	CONSTANT L : STD_LOGIC_VECTOR( 6 DOWNTO 0 ) := "1110001"; -- L
	CONSTANT A : STD_LOGIC_VECTOR( 6 DOWNTO 0 ) := "0001000"; -- A
	CONSTANT C : STD_LOGIC_VECTOR( 6 DOWNTO 0 ) := "1011101"; -- "

	TYPE MEMORIA IS ARRAY ( 5 DOWNTO 0 ) OF STD_LOGIC_VECTOR(BUS_DATOS'RANGE);
	
	CONSTANT ROM : MEMORIA := ( C, H, O, L, A, C );

	SIGNAL DATO : STD_LOGIC_VECTOR( BITS_BUS_DATOS-1 DOWNTO 0 );

	BEGIN

	DATO <= ROM( CONV_INTEGER(DIRECCION) );

	PBUF : PROCESS( CS, DATO )
	BEGIN
		IF ( CS = '1' ) THEN
			BUS_DATOS <= DATO;
		ELSE
			BUS_DATOS <= ( OTHERS => 'Z' );
		END IF;
	END PROCESS PBUF;

END MEMORIA;
