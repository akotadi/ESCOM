LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;

ENTITY IMP_DIS IS
	PORT(
		CLK, CLR, EN : IN STD_LOGIC;
		Q : INOUT STD_LOGIC_VECTOR(8 DOWNTO 0)
	);

	ATTRIBUTE PIN_NUMBERS OF IMP_DIS : ENTITY IS 
		"CLK:1 "		&
		"EN:2 "			&
		"CLR:13 "		&
		"Q(0):15 "		&
		"Q(1):16 "		&
		"Q(2):17 "		&
		"Q(3):18 "		&
		"Q(4):19 "		&
		"Q(5):20 "		&
		"Q(6):21";
END IMP_DIS;

ARCHITECTURE PRACTICA OF IMP_DIS IS

	CONSTANT Symbold : STD_LOGIC_VECTOR(6 DOWNTO 0) := "1000010";
	CONSTANT SymbolI : STD_LOGIC_VECTOR(6 DOWNTO 0) := "1001111";
	CONSTANT SymbolS : STD_LOGIC_VECTOR(6 DOWNTO 0) := "0100100";
	CONSTANT SymbolE : STD_LOGIC_VECTOR(6 DOWNTO 0) := "0110000";
	CONSTANT Symboln : STD_LOGIC_VECTOR(6 DOWNTO 0) := "0101010";
	CONSTANT SymbolO : STD_LOGIC_VECTOR(6 DOWNTO 0) := "0000001";
	CONSTANT Symbolg : STD_LOGIC_VECTOR(6 DOWNTO 0) := "0000100";
	CONSTANT Symbolt : STD_LOGIC_VECTOR(6 DOWNTO 0) := "1110000";
	CONSTANT SymbolA : STD_LOGIC_VECTOR(6 DOWNTO 0) := "0001000";
	CONSTANT SymbolL : STD_LOGIC_VECTOR(6 DOWNTO 0) := "1110001";

	CONSTANT Label00 : STD_LOGIC_VECTOR(1 DOWNTO 0) := "00";
	CONSTANT Label01 : STD_LOGIC_VECTOR(1 DOWNTO 0) := "01";
	CONSTANT Label10 : STD_LOGIC_VECTOR(1 DOWNTO 0) := "10";
	CONSTANT Label11 : STD_LOGIC_VECTOR(1 DOWNTO 0) := "11";

	CONSTANT q0 : STD_LOGIC_VECTOR(8 DOWNTO 0) := Label00&Symbold;
	CONSTANT q1 : STD_LOGIC_VECTOR(8 DOWNTO 0) := Label00&SymbolI;
	CONSTANT q2 : STD_LOGIC_VECTOR(8 DOWNTO 0) := Label00&SymbolS;
	CONSTANT q3 : STD_LOGIC_VECTOR(8 DOWNTO 0) := Label00&SymbolE;
	CONSTANT q4 : STD_LOGIC_VECTOR(8 DOWNTO 0) := Label00&Symboln;
	CONSTANT q5 : STD_LOGIC_VECTOR(8 DOWNTO 0) := Label00&SymbolO;
	CONSTANT q6 : STD_LOGIC_VECTOR(8 DOWNTO 0) := Label01&Symbold;
	CONSTANT q7 : STD_LOGIC_VECTOR(8 DOWNTO 0) := Label01&SymbolI;
	CONSTANT q8 : STD_LOGIC_VECTOR(8 DOWNTO 0) := Label00&Symbolg;
	CONSTANT q9 : STD_LOGIC_VECTOR(8 DOWNTO 0) := Label10&SymbolI;
	CONSTANT q10 : STD_LOGIC_VECTOR(8 DOWNTO 0) := Label00&Symbolt;
	CONSTANT q11 : STD_LOGIC_VECTOR(8 DOWNTO 0) := Label00&SymbolA;
	CONSTANT q12 : STD_LOGIC_VECTOR(8 DOWNTO 0) := Label00&SymbolL;

	BEGIN

		PROCESS(CLK, CLR)
			BEGIN
				IF (CLR = '1') THEN
					Q <= q0;
				ELSIF RISING_EDGE(CLK) THEN
					IF (EN = '1') THEN
						CASE Q IS
							WHEN q0 => Q <= q1;
							WHEN q1 => Q <= q2;
							WHEN q2 => Q <= q3;
							WHEN q3 => Q <= q4;
							WHEN q4 => Q <= q5;
							WHEN q5 => Q <= q6;
							WHEN q6 => Q <= q7;
							WHEN q7 => Q <= q8;
							WHEN q8 => Q <= q9;
							WHEN q9 => Q <= q10;
							WHEN q10 => Q <= q11;
							WHEN q11 => Q <= q12;
							WHEN OTHERS => Q <= q0;
						END CASE;
					END IF;
				END IF;
		END PROCESS;
END PRACTICA;