module variables ( 
	a,
	b,
	salida,
	cout
	) ;

input [3:0] a;
input [3:0] b;
inout [3:0] salida;
inout  cout;
