module suma ( 
	a,
	b,
	p
	) ;

input [1:0] a;
input [1:0] b;
inout [3:0] p;
