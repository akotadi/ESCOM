module suma ( 
	a,
	b,
	s,
	cout
	) ;

input [3:0] a;
input [3:0] b;
inout [3:0] s;
inout  cout;
