LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;

ENTITY ALARMAS IS

	PORT( 
		A,B,REF : in STD_LOGIC_VECTOR (2 downto 0);
		SEL: in STD_LOGIC;
		DISPLAY : out STD_LOGIC_VECTOR (6 downto 0)
	);

	ATTRIBUTE PIN_NUMBERS OF ALARMAS : ENTITY IS
		"DISPLAY(0):15 " &
		"DISPLAY(1):16 " &
		"DISPLAY(2):17 " &
		"DISPLAY(3):18 " &
		"DISPLAY(4):19 " &
		"DISPLAY(5):20 " &
		"DISPLAY(6):21";

END ALARMAS;

ARCHITECTURE CUADRO OF ALARMAS IS 

	SIGNAL SENSOR,CONDICION : STD_LOGIC_VECTOR(2 downto 0);
	
	BEGIN

		WITH SEL SELECT SENSOR <=
			A WHEN '0',
			B WHEN OTHERS;

		PCOMP : PROCESS(SENSOR,REF)
			BEGIN
				IF( SENSOR > REF ) THEN CONDICION <= "001";
				ELSIF( SENSOR = REF ) THEN CONDICION <= "010";
				ELSE CONDICION <= "100";
			END IF;
		END PROCESS PCOMP;

		DISPLAY <=
			"1111000" WHEN CONDICION = "001" ELSE
			"1001110" WHEN CONDICION = "100" ELSE
			"1001000";

END CUADRO;