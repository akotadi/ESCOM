LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_UNSIGNED.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

ENTITY CONTADOR IS 

	PORT( 
		CLK, CLR, LB, EB : IN STD_LOGIC;
		DB : IN STD_LOGIC_VECTOR(3 DOWNTO 0);
		B : INOUT STD_LOGIC_VECTOR(3 DOWNTO 0)
	);

END CONTADOR;



ARCHITECTURE PRACTICA OF CONTADOR IS 

	BEGIN

	CONT : PROCESS(CLK, CLR)

		BEGIN
			IF( CLR = '1' ) THEN
				B <= ( OTHERS => '0' );
			ELSIF RISING_EDGE(CLK) THEN
				IF ( LB = '1' ) THEN
					B <= DB;
				ELSIF ( EB = '1' ) THEN
					B <= B + 1;
				END IF;
			END IF;

	END PROCESS CONT;

END PRACTICA;