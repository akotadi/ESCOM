LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.ALL;

ENTITY program_memory IS
	GENERIC (
		BITS_BUS_DIR : INTEGER := 16;
		BITS_BUS_DATA : INTEGER := 25
	);

	Port ( 
		A : IN STD_LOGIC_VECTOR (BITS_BUS_DIR - 1 DOWNTO 0);
		D : IN STD_LOGIC_VECTOR (BITS_BUS_DATA - 1 DOWNTO 0)
	);
END program_memory;

ARCHITECTURE PROGRAMA OF program_memory IS

	-- CÓDIGOS DE OPERACIÓN
	CONSTANT OPCODE_TYPER : STD_LOGIC_VECTOR(4 DOWNTO 0) := "00000";
	CONSTANT OPCODE_LI : STD_LOGIC_VECTOR(4 DOWNTO 0) := "00001";
	CONSTANT OPCODE_LWI : STD_LOGIC_VECTOR(4 DOWNTO 0) := "00010";
	CONSTANT OPCODE_LW : STD_LOGIC_VECTOR(4 DOWNTO 0) := "10111";
	CONSTANT OPCODE_SWI : STD_LOGIC_VECTOR(4 DOWNTO 0) := "00011";
	CONSTANT OPCODE_SW : STD_LOGIC_VECTOR(4 DOWNTO 0) := "00100";
	CONSTANT OPCODE_ADDI : STD_LOGIC_VECTOR(4 DOWNTO 0) := "00101";
	CONSTANT OPCODE_SUBI : STD_LOGIC_VECTOR(4 DOWNTO 0) := "00110";
	CONSTANT OPCODE_ANDI : STD_LOGIC_VECTOR(4 DOWNTO 0) := "00111";
	CONSTANT OPCODE_ORI : STD_LOGIC_VECTOR(4 DOWNTO 0) := "01000";
	CONSTANT OPCODE_XORI : STD_LOGIC_VECTOR(4 DOWNTO 0) := "01001";
	CONSTANT OPCODE_NANDI : STD_LOGIC_VECTOR(4 DOWNTO 0) := "01010";
	CONSTANT OPCODE_NORI : STD_LOGIC_VECTOR(4 DOWNTO 0) := "01011";
	CONSTANT OPCODE_XNORI : STD_LOGIC_VECTOR(4 DOWNTO 0) := "01100";
	CONSTANT OPCODE_BEQI : STD_LOGIC_VECTOR(4 DOWNTO 0) := "01101";
	CONSTANT OPCODE_BNEI : STD_LOGIC_VECTOR(4 DOWNTO 0) := "01110";
	CONSTANT OPCODE_BLTI : STD_LOGIC_VECTOR(4 DOWNTO 0) := "01111";
	CONSTANT OPCODE_BLETI : STD_LOGIC_VECTOR(4 DOWNTO 0) := "10000";
	CONSTANT OPCODE_BGTI : STD_LOGIC_VECTOR(4 DOWNTO 0) := "10001";
	CONSTANT OPCODE_BGETI : STD_LOGIC_VECTOR(4 DOWNTO 0) := "10010";
	CONSTANT OPCODE_B : STD_LOGIC_VECTOR(4 DOWNTO 0) := "10011";
	CONSTANT OPCODE_CALL : STD_LOGIC_VECTOR(4 DOWNTO 0) := "10100";
	CONSTANT OPCODE_RET : STD_LOGIC_VECTOR(4 DOWNTO 0) := "10101";
	CONSTANT OPCODE_NOP : STD_LOGIC_VECTOR(4 DOWNTO 0) := "10110";

	-- CÓDIGOS DE FUNCIÓN
	CONSTANT FUNCODE_ADD : STD_LOGIC_VECTOR(3 DOWNTO 0) := X"0";
	CONSTANT FUNCODE_SUB : STD_LOGIC_VECTOR(3 DOWNTO 0) := X"1";
	CONSTANT FUNCODE_AND : STD_LOGIC_VECTOR(3 DOWNTO 0) := X"2";
	CONSTANT FUNCODE_OR : STD_LOGIC_VECTOR(3 DOWNTO 0) := X"3";
	CONSTANT FUNCODE_XOR : STD_LOGIC_VECTOR(3 DOWNTO 0) := X"4";
	CONSTANT FUNCODE_NAND : STD_LOGIC_VECTOR(3 DOWNTO 0) := X"5";
	CONSTANT FUNCODE_NOR : STD_LOGIC_VECTOR(3 DOWNTO 0) := X"6";
	CONSTANT FUNCODE_XNOR : STD_LOGIC_VECTOR(3 DOWNTO 0) := X"7";
	CONSTANT FUNCODE_NOT : STD_LOGIC_VECTOR(3 DOWNTO 0) := X"8";
	CONSTANT FUNCODE_SLL : STD_LOGIC_VECTOR(3 DOWNTO 0) := X"9";
	CONSTANT FUNCODE_SRL : STD_LOGIC_VECTOR(3 DOWNTO 0) := X"A";

	-- REGISTROS
	CONSTANT R0 : STD_LOGIC_VECTOR(3 DOWNTO 0) := X"0";
	CONSTANT R1 : STD_LOGIC_VECTOR(3 DOWNTO 0) := X"1";
	CONSTANT R2 : STD_LOGIC_VECTOR(3 DOWNTO 0) := X"2";
	CONSTANT R3 : STD_LOGIC_VECTOR(3 DOWNTO 0) := X"3";
	CONSTANT R4 : STD_LOGIC_VECTOR(3 DOWNTO 0) := X"4";
	CONSTANT R5 : STD_LOGIC_VECTOR(3 DOWNTO 0) := X"5";
	CONSTANT R6 : STD_LOGIC_VECTOR(3 DOWNTO 0) := X"6";
	CONSTANT R7 : STD_LOGIC_VECTOR(3 DOWNTO 0) := X"7";
	CONSTANT R8 : STD_LOGIC_VECTOR(3 DOWNTO 0) := X"8";
	CONSTANT R9 : STD_LOGIC_VECTOR(3 DOWNTO 0) := X"9";
	CONSTANT R10 : STD_LOGIC_VECTOR(3 DOWNTO 0) := X"A";
	CONSTANT R11 : STD_LOGIC_VECTOR(3 DOWNTO 0) := X"B";
	CONSTANT R12 : STD_LOGIC_VECTOR(3 DOWNTO 0) := X"C";
	CONSTANT R13 : STD_LOGIC_VECTOR(3 DOWNTO 0) := X"D";
	CONSTANT R14 : STD_LOGIC_VECTOR(3 DOWNTO 0) := X"E";
	CONSTANT R15 : STD_LOGIC_VECTOR(3 DOWNTO 0) := X"F";

	-- CAMPO SIN USO
	CONSTANT WU : STD_LOGIC_VECTOR(3 DOWNTO 0) := X"0";

	TYPE MEMORIA IS ARRAY (0 TO 2**BITS_BUS_DIR - 1) OF STD_LOGIC_VECTOR(D'RANGE);

	CONSTANT MEMP : MEMORIA := (
			--"00001 0000 0000 0000 0000 0001", 
			OPCODE_LI & R0 & X"0001", -- LI R0, #1
			--"00001 0001 0000 0000 0000 0111", 
			OPCODE_LI & R1 & X"0007", -- LI R1, #7
			OPCODE_TYPER & R1 & R1 & R0 & WU & FUNCODE_ADD, -- ADD R1, R1, R0
			OPCODE_SWI & R1 & X"0005", -- SWI R1, 5
			OPCODE_B & WU & X"0002", -- B CICLO
			OTHERS => (OTHERS => '0')
		);

	BEGIN

END PROGRAMA;