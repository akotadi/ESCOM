LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;

ENTITY FFS IS

	PORT( 
		J, K, T, D, S, R : IN STD_LOGIC;
		CLK, CLR : IN STD_LOGIC;
		SEL : IN STD_LOGIC_VECTOR(1 DOWNTO 0);
		-- QJK : INOUT STD_LOGIC; -- PODEMOS ESPECIFICARLE TERMINAL A UNA SEÑAL DE ESTA MANERA
		DISPLAY : OUT STD_LOGIC_VECTOR(5 DOWNTO 0)
	);

	ATTRIBUTE PIN_NUMBERS OF FFS : ENTITY IS
		"CLK:1 "		&
		"J:2 "			&
		"K:3 "			&
		"T:4 "			&
		"S:5 "			&
		"R:6 "			&
		"D:7 "			&
		"SEL(0):8 "		&
		"SEL(1):9 "		&
		"CLR:13 " 		&
		-- "QJK:15 " 	&
		"DISPLAY(0):16 " &
		"DISPLAY(1):17 " &
		"DISPLAY(2):18 " &
		"DISPLAY(3):19 " &
		"DISPLAY(4):20 " &
		"DISPLAY(5):21";

END FFS;

ARCHITECTURE PRACTICA OF FFS IS

	SIGNAL QJK, QT, QD, QSR, Q : STD_LOGIC;

	CONSTANT Visual0 : STD_LOGIC_VECTOR(5 DOWNTO 0) := "000000";
	CONSTANT Visual1 : STD_LOGIC_VECTOR(5 DOWNTO 0) := "100111";

	BEGIN

		FFJK : PROCESS( CLK, CLR ) -- J Y K SON SÍNCRONAS, DEPENDEN DEL CONTROL, POR ELLO NO SE COLOCAN
		BEGIN
			IF( CLR = '1' ) THEN
				QJK <= '0';
			ELSIF( CLK'EVENT AND CLK = '1' ) THEN
				QJK <= (NOT K AND QJK) OR (J AND NOT QJK);
			END IF;
		END PROCESS FFJK;

		FFT : PROCESS(CLK, CLR)
		BEGIN
			IF( CLR = '1' ) THEN
				QT <= '0';
			ELSIF( CLK'EVENT AND CLK = '1' ) THEN
				QT <= T XOR QT;
			END IF;
		END PROCESS FFT;

		FFD : PROCESS(CLK, CLR)
		BEGIN
			IF( CLR = '1' ) THEN
				QD <= '0';
			ELSIF( CLK'EVENT AND CLK = '1' ) THEN
				QD <= D;
			END IF;
		END PROCESS FFD;

		FFSR : PROCESS(CLK, CLR)
		BEGIN
			IF( CLR = '1' ) THEN
				QSR <= '0';
			ELSIF( CLK'EVENT AND CLK = '1' ) THEN
				QSR <= S OR (QSR AND NOT R);
			END IF;
		END PROCESS FFSR;

	--	WITH SEL SELECT Q <=
	--		QJK WHEN '00',
	--		QT WHEN '01',
	--		QD WHEN '10',
	--		QSR WHEN OTHERS;

	--	PCOMP : PROCESS(SENSOR,REF)
	--		BEGIN
	--			IF( SENSOR > REF ) THEN CONDICION <= "001";
	--			ELSIF( SENSOR = REF ) THEN CONDICION <= "010";
	--			ELSE CONDICION <= "100";
	--		END IF;
	--	END PROCESS PCOMP;

		 Q <=
			QJK WHEN SEL = "00" ELSE
			QT WHEN SEL = "01" ELSE
			QD WHEN SEL = "10" ELSE
			QSR;

		DISPLAY <=
			"000000" WHEN ( Q = '0' ) ELSE
			"100111";

END PRACTICA;