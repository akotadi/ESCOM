LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.ALL;

ENTITY CON_DEC_SHOW IS 	

	PORT( 
		CLK, CLR : IN STD_LOGIC;
		UNI : IN STD_LOGIC_VECTOR(3 DOWNTO 0);
		DEC : IN STD_LOGIC_VECTOR(2 DOWNTO 0);
		AN : INOUT STD_LOGIC_VECTOR(2 DOWNTO 0);
		DIS : OUT STD_LOGIC_VECTOR(6 DOWNTO 0)
	);

	ATTRIBUTE PIN_NUMBERS OF CON_DEC_SHOW : ENTITY IS 
		"CLK:1 "		&
		"CLR:13 "		&
		"UNI(0):11 "	&
		"UNI(1):10 "	&
		"UNI(2):9 "		&
		"UNI(3):8 "		&
		"DEC(0):7 "		&
		"DEC(1):6 "		&
		"DEC(2):5 "		&
		"AN(0):14 "		&
		"AN(1):23 "		&
		"AN(2):22 "		&
		"DIS(0):15 "	&
		"DIS(1):16 "	&
		"DIS(2):17 "	&
		"DIS(3):18 "	&
		"DIS(4):19 "	&
		"DIS(5):20 "	&
		"DIS(6):21";

END CON_DEC_SHOW;



ARCHITECTURE PRACTICA OF CON_DEC_SHOW IS 

	CONSTANT Symbol0 : STD_LOGIC_VECTOR(6 DOWNTO 0) := "0000001";
	CONSTANT Symbol1 : STD_LOGIC_VECTOR(6 DOWNTO 0) := "1001111";
	CONSTANT Symbol2 : STD_LOGIC_VECTOR(6 DOWNTO 0) := "0010010";
	CONSTANT Symbol3 : STD_LOGIC_VECTOR(6 DOWNTO 0) := "0000110";
	CONSTANT Symbol4 : STD_LOGIC_VECTOR(6 DOWNTO 0) := "1001100";
	CONSTANT Symbol5 : STD_LOGIC_VECTOR(6 DOWNTO 0) := "0100100";
	CONSTANT Symbol6 : STD_LOGIC_VECTOR(6 DOWNTO 0) := "0100000";
	CONSTANT Symbol7 : STD_LOGIC_VECTOR(6 DOWNTO 0) := "0001111";
	CONSTANT Symbol8 : STD_LOGIC_VECTOR(6 DOWNTO 0) := "0000000";
	CONSTANT Symbol9 : STD_LOGIC_VECTOR(6 DOWNTO 0) := "0000100";

	CONSTANT BCD0 : STD_LOGIC_VECTOR(3 DOWNTO 0) := "0000";
	CONSTANT BCD1 : STD_LOGIC_VECTOR(3 DOWNTO 0) := "0001";
	CONSTANT BCD2 : STD_LOGIC_VECTOR(3 DOWNTO 0) := "0010";
	CONSTANT BCD3 : STD_LOGIC_VECTOR(3 DOWNTO 0) := "0011";
	CONSTANT BCD4 : STD_LOGIC_VECTOR(3 DOWNTO 0) := "0100";
	CONSTANT BCD5 : STD_LOGIC_VECTOR(3 DOWNTO 0) := "0101";
	CONSTANT BCD6 : STD_LOGIC_VECTOR(3 DOWNTO 0) := "0110";
	CONSTANT BCD7 : STD_LOGIC_VECTOR(3 DOWNTO 0) := "0111";
	CONSTANT BCD8 : STD_LOGIC_VECTOR(3 DOWNTO 0) := "1000";
	CONSTANT BCD9 : STD_LOGIC_VECTOR(3 DOWNTO 0) := "1001";

	SIGNAL BCD : STD_LOGIC_VECTOR(3 DOWNTO 0); 
--	SIGNAL CENT : STD_LOGIC_VECTOR(3 DOWNTO 0);

	BEGIN

--	CENT <= ( OTHERS => '0' );

	CONT_AN : PROCESS(CLK, CLR)
		BEGIN
			IF( CLR = '1' ) THEN
				AN <= "110";
			ELSIF RISING_EDGE(CLK) THEN
				AN <= TO_STDLOGICVECTOR( TO_BITVECTOR( AN ) ROL 1 );
			END IF;
	END PROCESS CONT_AN;

	MUX : PROCESS(AN, UNI, DEC)
		BEGIN
			CASE AN IS
				WHEN "110" => BCD <= UNI;
				WHEN "101" => 
					BCD <= '0'&DEC;
--					BCD(3) <= '0';
--					BCD(2) <= DEC(2);
--					BCD(1) <= DEC(1);
--					BCD(0) <= DEC(0);
				WHEN "011" => BCD <= (OTHERS => '0');
				WHEN OTHERS => BCD <= (OTHERS => '0');
			END CASE;
	END PROCESS MUX;

	DISPLAY : PROCESS(BCD)
		BEGIN
			CASE BCD IS
				WHEN BCD0 => DIS <= Symbol0;
				WHEN BCD1 => DIS <= Symbol1;
				WHEN BCD2 => DIS <= Symbol2;
				WHEN BCD3 => DIS <= Symbol3;
				WHEN BCD4 => DIS <= Symbol4;
				WHEN BCD5 => DIS <= Symbol5;
				WHEN BCD6 => DIS <= Symbol6;
				WHEN BCD7 => DIS <= Symbol7;
				WHEN BCD8 => DIS <= Symbol8;
				WHEN BCD9 => DIS <= Symbol9;
				WHEN OTHERS => DIS <= (OTHERS => '-');
			END CASE;
	END PROCESS DISPLAY;

END PRACTICA;