LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_UNSIGNED.ALL;

ENTITY MARQUESINA IS 

	GENERIC (
		BITS_BUS_DIR : INTEGER := 3;
		BITS_BUS_DATOS : INTEGER := 7
	);

	PORT(
		DIRECCION : IN STD_LOGIC_VECTOR( BITS_BUS_DIR-1 DOWNTO 0 );
		DIS : OUT STD_LOGIC_VECTOR( BITS_BUS_DATOS-1 DOWNTO 0 );
		AN : INOUT STD_LOGIC_VECTOR(2 DOWNTO 0);
		CLK, CLR : IN STD_LOGIC
	);

	ATTRIBUTE PIN_NUMBERS OF MARQUESINA : ENTITY IS 
		"CLK:1 "				&
		"CLR:13 "				&
		"DIRECCION(0):6 "		&
		"DIRECCION(1):5 "		&
		"DIRECCION(2):4 "		&
		"AN(0):14 "				&
		"AN(1):23 "				&
		"AN(2):22 "				&
		"DIS(0):15 "			&
		"DIS(1):16 "			&
		"DIS(2):17 "			&
		"DIS(3):18 "			&
		"DIS(4):19 "			&
		"DIS(5):20 "			&
		"DIS(6):21";

END MARQUESINA;

ARCHITECTURE PRACTICA OF MARQUESINA IS 

	CONSTANT Symbold : STD_LOGIC_VECTOR(6 DOWNTO 0) := "1000010"; -- 42
	CONSTANT SymbolI : STD_LOGIC_VECTOR(6 DOWNTO 0) := "1001111"; -- 4F
	CONSTANT SymbolS : STD_LOGIC_VECTOR(6 DOWNTO 0) := "0100100"; -- 24
	CONSTANT SymbolE : STD_LOGIC_VECTOR(6 DOWNTO 0) := "0110000"; -- 30
	CONSTANT Symboln : STD_LOGIC_VECTOR(6 DOWNTO 0) := "0101010"; -- 2C
	CONSTANT SymbolO : STD_LOGIC_VECTOR(6 DOWNTO 0) := "0000001"; -- 01
	CONSTANT Symbolc : STD_LOGIC_VECTOR(6 DOWNTO 0) := "1110111"; -- 77

	TYPE MEMORIA IS ARRAY ( 7 DOWNTO 0 ) OF STD_LOGIC_VECTOR( BITS_BUS_DATOS-1 DOWNTO 0 );
	
	CONSTANT ROM2 : MEMORIA := ( SymbolO, Symboln, SymbolE, SymbolS, SymbolI, Symbold, Symbolc, Symbolc );
	CONSTANT ROM1 : MEMORIA := ( Symbolc, SymbolO, Symboln, SymbolE, SymbolS, SymbolI, Symbold, Symbolc );
	CONSTANT ROM0 : MEMORIA := ( Symbolc, Symbolc, SymbolO, Symboln, SymbolE, SymbolS, SymbolI, Symbold );

	SIGNAL DISP2 : STD_LOGIC_VECTOR( BITS_BUS_DATOS-1 DOWNTO 0 );
	SIGNAL DISP1 : STD_LOGIC_VECTOR( BITS_BUS_DATOS-1 DOWNTO 0 );
	SIGNAL DISP0 : STD_LOGIC_VECTOR( BITS_BUS_DATOS-1 DOWNTO 0 );

	BEGIN

	CONT_AN : PROCESS( CLK, CLR )
		BEGIN
			IF( CLR = '1' ) THEN
				AN <= "110";
			ELSIF RISING_EDGE(CLK) THEN
				AN <= TO_STDLOGICVECTOR( TO_BITVECTOR( AN ) ROL 1 );
			END IF;
	END PROCESS CONT_AN;

	DISP2 <= ROM2( CONV_INTEGER(DIRECCION) );

	DISP1 <= ROM1( CONV_INTEGER(DIRECCION) );

	DISP0 <= ROM0( CONV_INTEGER(DIRECCION) );

	MUX : PROCESS( AN, DISP0, DISP1, DISP2 )
		BEGIN
			CASE AN IS
				WHEN "110" => DIS <= DISP0;
				WHEN "101" => DIS <= DISP1;
				WHEN "011" => DIS <= DISP2;
				WHEN OTHERS => DIS <= ( OTHERS => '-' );
			END CASE;
	END PROCESS MUX;

END PRACTICA;
