LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_UNSIGNED.ALL;

ENTITY MARQUESINA IS 

	GENERIC (
		BITS_BUS_DIR : INTEGER := 4;
		BITS_BUS_DATOS : INTEGER := 7
	);

	PORT(
		VENTANA : IN STD_LOGIC_VECTOR( 2 DOWNTO 0 );
		DIS : OUT STD_LOGIC_VECTOR( 6 DOWNTO 0 );
		AN : INOUT STD_LOGIC_VECTOR(2 DOWNTO 0);
		CLK, CLR : IN STD_LOGIC
	);

	ATTRIBUTE PIN_NUMBERS OF MARQUESINA : ENTITY IS 
		"CLK:1 "				&
		"CLR:13 "				&
		"VENTANA(0):6 "			&
		"VENTANA(1):5 "			&
		"VENTANA(2):4 "			&
		"AN(0):14 "				&
		"AN(1):23 "				&
		"AN(2):22 "				&
		"DIS(0):15 "			&
		"DIS(1):16 "			&
		"DIS(2):17 "			&
		"DIS(3):18 "			&
		"DIS(4):19 "			&
		"DIS(5):20 "			&
		"DIS(6):21";

END MARQUESINA;

ARCHITECTURE PRACTICA OF MARQUESINA IS 

	CONSTANT SymbolE : STD_LOGIC_VECTOR(6 DOWNTO 0) := "0110000"; -- 30
	CONSTANT SymbolS : STD_LOGIC_VECTOR(6 DOWNTO 0) := "0100100"; -- 24
	CONSTANT SymbolC : STD_LOGIC_VECTOR(6 DOWNTO 0) := "0110001"; -- 31
	CONSTANT SymbolO : STD_LOGIC_VECTOR(6 DOWNTO 0) := "0000001"; -- 01
	CONSTANT Symboln : STD_LOGIC_VECTOR(6 DOWNTO 0) := "0101010"; -- 2A
	CONSTANT SymbolX : STD_LOGIC_VECTOR(6 DOWNTO 0) := "1110111"; -- 77

	TYPE MEMORIA IS ARRAY ( 9 DOWNTO 0 ) OF STD_LOGIC_VECTOR( BITS_BUS_DATOS-1 DOWNTO 0 );
	
	CONSTANT ROM : MEMORIA := ( SymbolX, SymbolX, Symboln, Symboln, SymbolO, SymbolC, SymbolS, SymbolE, SymbolX, SymbolX );

	SIGNAL DATOS : STD_LOGIC_VECTOR( BITS_BUS_DATOS-1 DOWNTO 0 );

	SIGNAL DESP : STD_LOGIC_VECTOR( 2 DOWNTO 0 );

	BEGIN

	CONT_AN : PROCESS( CLK, CLR )
		BEGIN
			IF( CLR = '1' ) THEN
				AN <= "110";
			ELSIF RISING_EDGE(CLK) THEN
				AN <= TO_STDLOGICVECTOR( TO_BITVECTOR( AN ) ROL 1 );
			END IF;
	END PROCESS CONT_AN;

	-- Añadir suma con ecuaciones

	SUMADOR : PROCESS (VENTANA, DESP)
		BEGIN

	END PROCESS SUMADOR;

	DIS <= ROM( CONV_INTEGER(VENTANA) + CONV_INTEGER(DESP) );

	CONV_COD : PROCESS( AN )
		BEGIN
			CASE AN IS
				WHEN "110" => DESP <= "010";
				WHEN "101" => DESP <= "001";
				WHEN "011" => DESP <= "000";
				WHEN OTHERS => DESP <= ( OTHERS => '-' );
			END CASE;
	END PROCESS CONV_COD;

END PRACTICA;
