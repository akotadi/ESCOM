module compuertas ( 
	a1,
	a2,
	a3,
	a4,
	b1,
	b2,
	b3,
	b4,
	sel,
	cout,
	s1,
	s2,
	s3,
	s4
	) ;

input  a1;
input  a2;
input  a3;
input  a4;
input  b1;
input  b2;
input  b3;
input  b4;
input  sel;
inout  cout;
inout  s1;
inout  s2;
inout  s3;
inout  s4;
