LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.ALL;

ENTITY COMPUERTAS IS
	PORT(
			AMS: in STD_LOGIC;
			BMS: in STD_LOGIC;
			CinSC: in STD_LOGIC;
			CoSC: out STD_LOGIC;
			CMS: out STD_LOGIC;
			SSC: out STD_LOGIC;
			SMS: out STD_LOGIC;
			AMR: in STD_LOGIC;
			BMR: in STD_LOGIC;
			PiRC: in STD_LOGIC;
			RMR: out STD_LOGIC;
			PMR: out STD_LOGIC;
			PoRC: out STD_LOGIC;
			RRC: out STD_LOGIC
		);

	ATTRIBUTE PIN_NUMBERS OF COMPUERTAS: ENTITY IS
	"AMS:1 BMS:2 CinSC:3 AMR:4 BMR:5 PiRC:6"
	& " SMS:14 CMS:15 CoSC:16 SSC:17"
	& " RMR:18 PMR:19 PoRC:20 RRC:21";

END COMPUERTAS;

ARCHITECTURE BEHAVIORAL OF COMPUERTAS IS
	BEGIN
		SMS<= AMS XOR BMS;
		CMS<= AMS AND BMS;
		CoSC<= ((AMS XOR BMS)AND CinSC) OR (AMS AND BMS);
		SSC<= (AMS XOR BMS) XOR CinSC;

		RMR<= AMR XOR BMR;
		PMR<= NOT(AMR) AND BMR;
		RRC<= (BMR XOR PiRC) XOR AMR;
		PoRC<= (NOT(AMR) AND PiRC) OR (NOT(AMR) AND BMR) OR (BMR AND PiRC);

	END BEHAVIORAL;
