LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_UNSIGNED.ALL;

ENTITY MARQUESINA IS 

	GENERIC (
		BITS_BUS_DIR : INTEGER := 4;
		BITS_BUS_DATOS : INTEGER := 4
	);

	PORT(
		DIRECCION : IN STD_LOGIC_VECTOR( BITS_BUS_DIR-1 DOWNTO 0 );
		DIS : OUT STD_LOGIC_VECTOR( 6 DOWNTO 0 );
		AN : INOUT STD_LOGIC_VECTOR(2 DOWNTO 0);
		CLK, CLR : IN STD_LOGIC
	);

	ATTRIBUTE PIN_NUMBERS OF MARQUESINA : ENTITY IS 
		"CLK:1 "				&
		"CLR:13 "				&
		"DIRECCION(0):7 "		&
		"DIRECCION(1):6 "		&
		"DIRECCION(2):5 "		&
		"DIRECCION(3):4 "		&
		"AN(0):14 "				&
		"AN(1):23 "				&
		"AN(2):22 "				&
		"DIS(0):15 "			&
		"DIS(1):16 "			&
		"DIS(2):17 "			&
		"DIS(3):18 "			&
		"DIS(4):19 "			&
		"DIS(5):20 "			&
		"DIS(6):21";

END MARQUESINA;

ARCHITECTURE PRACTICA OF MARQUESINA IS 

	CONSTANT Symbold : STD_LOGIC_VECTOR(6 DOWNTO 0) := "1000010"; -- 42
	CONSTANT SymbolI : STD_LOGIC_VECTOR(6 DOWNTO 0) := "1001111"; -- 4F
	CONSTANT SymbolS : STD_LOGIC_VECTOR(6 DOWNTO 0) := "0100100"; -- 24
	CONSTANT SymbolE : STD_LOGIC_VECTOR(6 DOWNTO 0) := "0110000"; -- 30
	CONSTANT Symboln : STD_LOGIC_VECTOR(6 DOWNTO 0) := "0101010"; -- 2A
	CONSTANT SymbolO : STD_LOGIC_VECTOR(6 DOWNTO 0) := "0000001"; -- 01
	CONSTANT Symbolc : STD_LOGIC_VECTOR(6 DOWNTO 0) := "1110111"; -- 77
	CONSTANT Symbolg : STD_LOGIC_VECTOR(6 DOWNTO 0) := "0000100"; -- 04
	CONSTANT Symbolt : STD_LOGIC_VECTOR(6 DOWNTO 0) := "1110000"; -- 70
	CONSTANT SymbolA : STD_LOGIC_VECTOR(6 DOWNTO 0) := "0001000"; -- 08
	CONSTANT SymbolL : STD_LOGIC_VECTOR(6 DOWNTO 0) := "1110001"; -- 71

	CONSTANT Codc : STD_LOGIC_VECTOR(3 DOWNTO 0) := "0000"; -- 0
	CONSTANT Codd : STD_LOGIC_VECTOR(3 DOWNTO 0) := "0001"; -- 1
	CONSTANT CodI : STD_LOGIC_VECTOR(3 DOWNTO 0) := "0011"; -- 3
	CONSTANT CodS : STD_LOGIC_VECTOR(3 DOWNTO 0) := "0010"; -- 2
	CONSTANT CodE : STD_LOGIC_VECTOR(3 DOWNTO 0) := "0110"; -- 6
	CONSTANT Codn : STD_LOGIC_VECTOR(3 DOWNTO 0) := "0111"; -- 7
	CONSTANT CodO : STD_LOGIC_VECTOR(3 DOWNTO 0) := "0101"; -- 5
	CONSTANT Codg : STD_LOGIC_VECTOR(3 DOWNTO 0) := "0100"; -- 4
	CONSTANT Codt : STD_LOGIC_VECTOR(3 DOWNTO 0) := "1100"; -- C
	CONSTANT CodA : STD_LOGIC_VECTOR(3 DOWNTO 0) := "1101"; -- D
	CONSTANT CodL : STD_LOGIC_VECTOR(3 DOWNTO 0) := "1111"; -- F
	CONSTANT CodX : STD_LOGIC_VECTOR(3 DOWNTO 0) := "1110"; -- E

	TYPE MEMORIA IS ARRAY ( 15 DOWNTO 0 ) OF STD_LOGIC_VECTOR( BITS_BUS_DATOS-1 DOWNTO 0 );
	
	CONSTANT ROM2 : MEMORIA := ( CodL, CodA, Codt, CodI, Codg, CodI, Codd, Codc, CodO, Codn, CodE, CodS, CodI, Codd, Codc, Codc );
	CONSTANT ROM1 : MEMORIA := ( Codc, CodL, CodA, Codt, CodI, Codg, CodI, Codd, Codc, CodO, Codn, CodE, CodS, CodI, Codd, Codc );
	CONSTANT ROM0 : MEMORIA := ( Codc, Codc, CodL, CodA, Codt, CodI, Codg, CodI, Codd, Codc, CodO, Codn, CodE, CodS, CodI, Codd );

	SIGNAL DISP2 : STD_LOGIC_VECTOR( BITS_BUS_DATOS-1 DOWNTO 0 );
	SIGNAL DISP1 : STD_LOGIC_VECTOR( BITS_BUS_DATOS-1 DOWNTO 0 );
	SIGNAL DISP0 : STD_LOGIC_VECTOR( BITS_BUS_DATOS-1 DOWNTO 0 );

	SIGNAL COD_DIS : STD_LOGIC_VECTOR( 3 DOWNTO 0 );

	BEGIN

	CONT_AN : PROCESS( CLK, CLR )
		BEGIN
			IF( CLR = '1' ) THEN
				AN <= "110";
			ELSIF RISING_EDGE(CLK) THEN
				AN <= TO_STDLOGICVECTOR( TO_BITVECTOR( AN ) ROL 1 );
			END IF;
	END PROCESS CONT_AN;

	DISP2 <= ROM2( CONV_INTEGER(DIRECCION) );

	DISP1 <= ROM1( CONV_INTEGER(DIRECCION) );

	DISP0 <= ROM0( CONV_INTEGER(DIRECCION) );

	MUX : PROCESS( AN )
		BEGIN
			CASE AN IS
				WHEN "110" => COD_DIS <= DISP0;
				WHEN "101" => COD_DIS <= DISP1;
				WHEN "011" => COD_DIS <= DISP2;
				WHEN OTHERS => COD_DIS <= CodX;
			END CASE;
	END PROCESS MUX;

	CONV_COD : PROCESS( COD_DIS )
		BEGIN
			CASE COD_DIS IS
				WHEN Codc => DIS <= Symbolc;
				WHEN Codd => DIS <= Symbold;
				WHEN CodI => DIS <= SymbolI;
				WHEN CodS => DIS <= SymbolS;
				WHEN CodE => DIS <= SymbolE;
				WHEN Codn => DIS <= Symboln;
				WHEN CodO => DIS <= SymbolO;
				WHEN Codg => DIS <= Symbolg;
				WHEN Codt => DIS <= Symbolt;
				WHEN CodA => DIS <= SymbolA;
				WHEN CodL => DIS <= SymbolL;
				WHEN OTHERS => DIS <= ( OTHERS => '-' );
			END CASE;
	END PROCESS CONV_COD;

END PRACTICA;
