module variables ( 
	a,
	b,
	c,
	d,
	c0,
	c1,
	a1,
	c2,
	b1,
	c11,
	d1
	) ;

input  a;
input  b;
input  c;
input  d;
inout  c0;
inout  c1;
inout  a1;
inout  c2;
inout  b1;
inout  c11;
inout  d1;
