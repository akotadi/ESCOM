LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_UNSIGNED.ALL;

ENTITY ROM IS 

	GENERIC (
		BITS_BUS_DIR : INTEGER := 7;
		BITS_BUS_DATOS : INTEGER := 8
	);

	PORT(
		DIRECCION : IN STD_LOGIC_VECTOR( BITS_BUS_DIR-1 DOWNTO 0 );
		BUS_DATOS : OUT STD_LOGIC_VECTOR( BITS_BUS_DATOS-1 DOWNTO 0 );
		CS : IN STD_LOGIC
	);

END ROM;

ARCHITECTURE MEMORIA OF ROM IS 

	TYPE MEMORIA IS ARRAY ( 0 TO 2**BITS_BUS_DIR-1 ) OF STD_LOGIC_VECTOR(BUS_DATOS'RANGE);
	
	CONSTANT ROM : MEMORIA := ( 
		X"03",
		X"45",
		X"A3",
		X"B2",
		OTHERS => X"00"
	);

	SIGNAL DATO : STD_LOGIC_VECTOR( BITS_BUS_DATOS-1 DOWNTO 0 );

	BEGIN

	DATO <= ROM( CONV_INTEGER(DIRECCION) );

	PBUF : PROCESS( CS, DATO )
	BEGIN
		IF ( CS = '1' ) THEN
			BUS_DATOS <= DATO;
		ELSE
			BUS_DATOS <= ( OTHERS => 'Z' );
		END IF;
	END PROCESS PBUF;

END MEMORIA;
