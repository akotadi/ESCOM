LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.ALL;

ENTITY DECO IS
	PORT(
		E	:IN STD_LOGIC_VECTOR(2 DOWNTO 0);
	DISPLAY	:OUT STD_LOGIC_VECTOR(6 DOWNTO 0)
		);
END DECO;

ARCHITECTURE ADECO OF DECO IS
BEGIN
	PDECO : PROCESS( E )
	BEGIN
			CASE E IS
					WHEN "000" => DISPLAY <= "0000000"; --8
					WHEN "001" => DISPLAY <= "000110"; --9
					WHEN "010" => DISPLAY <= "010010"; --5
					WHEN "011" => DISPLAY <= "010000"; --6
					WHEN "100" => DISPLAY <= "000001"; --0
					WHEN "101" => DISPLAY <= "101111"; --1
					WHEN "110" => DISPLAY <= "001111"; --7
					WHEN OTHERS => DISPLAY <= "0011000"; --1
			 END CASE;
	END PROCESS PDECO;
END ADECO;
