LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;

ENTITY CONTADOR IS 

	GENERIC( 
		N : INTEGER := 7 
	);

	PORT( 
		CLK, CLR: IN STD_LOGIC;
		F : IN STD_LOGIC_VECTOR(3 DOWNTO 0);
		C : INOUT STD_LOGIC_VECTOR(2 DOWNTO 0);
		DIS : INOUT STD_LOGIC_VECTOR(N-1 DOWNTO 0)
	);

	ATTRIBUTE PIN_NUMBERS OF CONTADOR : ENTITY IS 
		"CLK:1 "			&
		"F(0):8 "			&
		"F(1):9 "			&
		"F(2):10 "			&
		"F(3):11 "			&
		"C(0):14 "			&
		"C(1):22 "			&
		"C(2):23 "			&
		"DIS(0):15 "		&
		"DIS(1):16 "		&
		"DIS(2):17 "		&
		"DIS(3):18 "		&
		"DIS(4):19 "		&
		"DIS(5):20 "		&
		"DIS(6):21 "		&
		"CLR:13";

END CONTADOR;



ARCHITECTURE PRACTICA OF CONTADOR IS 

	SIGNAL L : STD_LOGIC;
	SIGNAL BUTTON : STD_LOGIC_VECTOR(6 DOWNTO 0);

	CONSTANT Symbol0 : STD_LOGIC_VECTOR(6 DOWNTO 0) := "0000001";
	CONSTANT Symbol1 : STD_LOGIC_VECTOR(6 DOWNTO 0) := "1001111";
	CONSTANT Symbol2 : STD_LOGIC_VECTOR(6 DOWNTO 0) := "0010010";
	CONSTANT Symbol3 : STD_LOGIC_VECTOR(6 DOWNTO 0) := "0000110";
	CONSTANT Symbol4 : STD_LOGIC_VECTOR(6 DOWNTO 0) := "1001100";
	CONSTANT Symbol5 : STD_LOGIC_VECTOR(6 DOWNTO 0) := "0100100";
	CONSTANT Symbol6 : STD_LOGIC_VECTOR(6 DOWNTO 0) := "0100000";
	CONSTANT Symbol7 : STD_LOGIC_VECTOR(6 DOWNTO 0) := "0001111";
	CONSTANT Symbol8 : STD_LOGIC_VECTOR(6 DOWNTO 0) := "0000000";
	CONSTANT Symbol9 : STD_LOGIC_VECTOR(6 DOWNTO 0) := "0001100";
	CONSTANT SymbolA : STD_LOGIC_VECTOR(6 DOWNTO 0) := "0001000";
	CONSTANT Symbolg : STD_LOGIC_VECTOR(6 DOWNTO 0) := "0000100";

	BEGIN

	L <= NOT ( F(0) AND F(1) AND F(2) AND F(3) );

	CONT_AN : PROCESS(CLK, CLR)
		BEGIN
			IF( CLR = '1' ) THEN
				C <= "110";

			ELSIF RISING_EDGE(CLK) THEN
				C <= TO_STDLOGICVECTOR( TO_BITVECTOR( C ) ROL 1 );
			END IF;
	END PROCESS CONT_AN;

	DISPLAY : PROCESS(F, C)
		BEGIN
			CASE F&C IS
				WHEN "1110011" => BUTTON <= Symbol1;
				WHEN "1101011" => BUTTON <= Symbol4;
				WHEN "1011011" => BUTTON <= Symbol7;
				WHEN "0111011" => BUTTON <= SymbolA;
				WHEN "1110101" => BUTTON <= Symbol2;
				WHEN "1101101" => BUTTON <= Symbol5;
				WHEN "1011101" => BUTTON <= Symbol8;
				WHEN "0111101" => BUTTON <= Symbol0;
				WHEN "1110110" => BUTTON <= Symbol3;
				WHEN "1101110" => BUTTON <= Symbol6;
				WHEN "1011110" => BUTTON <= Symbol9;
				WHEN "0111110" => BUTTON <= Symbolg;
				WHEN OTHERS => BUTTON <= ( OTHERS => '-' );
			END CASE;
	END PROCESS DISPLAY;

	REG : PROCESS(CLK, CLR)
		BEGIN
			IF ( CLR = '1' ) THEN
				DIS <= (OTHERS => '1');
			ELSIF RISING_EDGE(CLK) THEN
				IF ( L = '1' ) THEN
					DIS <= BUTTON;
				ELSE
					DIS <= DIS;
				END IF;
			END IF;
	END PROCESS REG;

END PRACTICA;