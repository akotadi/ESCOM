LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.ALL;

ENTITY SUMA IS
	PORT(
		A,B: in STD_LOGIC_VECTOR(1 downto 0);
		P: out STD_LOGIC_VECTOR(3 downto 0)
		);

  
	ATTRIBUTE PIN_NUMBERS OF SUMA: ENTITY IS
	"P(0):18 P(1):17 P(2):16 P(3):15";
END SUMA;

ARCHITECTURE BEHAVIORAL OF SUMA IS
begin
	P(0)<=A(0)AND B(0);
	P(1)<=(A(1) AND B(0)) XOR (A(0) AND B(1));
	P(2)<=(A(1) AND B(1)) XOR ((A(1) AND B(0)) AND (A(0) AND B(1)));
	P(3)<=(A(1) AND B(1)) AND ((A(1) AND B(0)) AND (A(0) AND B(1)));

	END BEHAVIORAL;